library ieee;
use     ieee.std_logic_1164.all;

package utilities is
  
	type ball_direction_h_type is (left, right);
	type ball_direction_v_type is (up, down);
  
end package;